module fetch_controller (
    input [6:0] opcode,
    output ex_signals,
    output mem_signals,
    output wb_signals
);


endmodule