module fetch_controller (
    input [6:0] opcode;
)


endmodule