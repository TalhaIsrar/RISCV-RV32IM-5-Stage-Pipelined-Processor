module rv32i_core(
    input clk,
    input rst
);

endmodule