// OPCODES
`define OPCODE_RTYPE 7'b0110011