module pc(

)


endmodule